/*                                                                      
    Designer   : Renyangang               
                                                                            
    Licensed under the Apache License, Version 2.0 (the "License");         
    you may not use this file except in compliance with the License.        
    You may obtain a copy of the License at                                 
                                                                            
        http://www.apache.org/licenses/LICENSE-2.0                          
                                                                            
    Unless required by applicable law or agreed to in writing, software    
    distributed under the License is distributed on an "AS IS" BASIS,       
    WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
    See the License for the specific language governing permissions and     
    limitations under the License. 
*/
module t(
    input clk,
    input rst,
    output reg [3:0] leds
);

    always @(posedge clk or rst) begin
        if (!rst) begin
            leds <= 4'b0001;
        end
        else begin
            leds <= {leds[2:0], leds[3]};
        end
    end
endmodule